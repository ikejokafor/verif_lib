`ifndef	__VERIFICATION_DEFS__
`define	__VERIFICATION_DEFS__


typedef enum bit {TRUE = 1, FALSE = 0} bool;
typedef bit [127:0] mem_queue_64_t[$];


`endif